
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

-- 实体 AC_A 寄存器
ENTITY AC_A IS
PORT(
     LOAD_A 	: IN 	STD_LOGIC;
	  clk 		: IN 	STD_LOGIC;
	  Data_in 	: IN 	STD_LOGIC_VECTOR(15 DOWNTO 0);
	  A 			: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
);
END AC_A;

-- 结构体 func
ARCHITECTURE accu OF AC_A IS
	-- 变量声明 func

-- 功能 func
BEGIN
	PROCESS(clk,LOAD_A,data_in)	-- 进程 变量输入
	BEGIN
		IF clk'event AND clk = '1' THEN
			IF LOAD_A = '1' THEN
				A <= Data_in;
			END IF;
		END IF;
	END PROCESS;
END accu; -- 结构体 结束
	  

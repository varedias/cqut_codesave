LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY SAVER IS
PORT(
    Data_in   : IN    STD_LOGIC_VECTOR(15 DOWNTO 0);
    A         : OUT   STD_LOGIC_VECTOR(15 DOWNTO 0)
  
);
END SAVER;

ARCHITECTURE accu OF SAVER IS
BEGIN
    PROCESS (Data_in) 
    BEGIN
            A <= Data_in; 
      
        
    END PROCESS;
END accu;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PC IS
PORT(
	clk 			: IN 		STD_LOGIC;	
	Reset 		: IN 		STD_LOGIC;	
	LOAD_PC 		: IN 		STD_LOGIC;	
	INCR_PC 		: IN 		STD_LOGIC;	
	Addr_in	: IN		STD_LOGIC_VECTOR(7 DOWNTO 0);	
	PC_out 		: INOUT 	STD_LOGIC_VECTOR(7 DOWNTO 0)	
);
END PC;


ARCHITECTURE BEHAVE OF PC IS


BEGIN
	PROCESS(CLK,Reset,LOAD_PC,INCR_PC)	
	BEGIN
		IF Reset = '1' THEN
			PC_out <= X"00";
		ELSIF clk'event AND clk = '1' THEN
			IF LOAD_PC = '0' AND INCR_PC = '1' THEN		
				PC_out <=PC_out+X"01";
		   ELSIF LOAD_PC = '1' AND INCR_PC = '0' THEN	
		      PC_out <= Addr_in;
		   END IF;
		END IF;
	END PROCESS;
END BEHAVE; 
		  